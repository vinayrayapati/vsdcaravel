module scl_decap_12 ();
    // Voltage supply signals
    supply1 VPWR;
    supply0 VGND;
    supply1 VPB ;
    supply0 VNB ;

    scl_decap base ();

endmodule

module scl_decap ();
     // No contents.
endmodule
